/**
	\author: 	Trasier
	\date: 		2017/5/10
	\brief: 	TOY of the Controller
*/
module toyCU (

);

endmodule
