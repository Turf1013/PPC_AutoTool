/*
 * Description: This module is all about definition of default.
 * Author: ZengYX
 * Date:   2014.8.7
 */
 
`define MUX_D_DEFAULT	0 